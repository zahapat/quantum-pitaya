package generics is

    constant INT_BYPASS_DSP : integer := 0;
    constant INT_WHOLE_DDC_LOCOSC_OUT_FREQ_MHZ : integer := 25;
    constant INT_DECIMAL_DDC_LOCOSC_OUT_FREQ_MHZ : integer := 0;
    constant INT_DDC_NUMBER_OF_TAPS : integer := 15;
    constant INT_DDC_COEF_WIDTH : integer := 15;
    constant INT_DDC_OUT_DATA_WIDTH : integer := 20;
    constant INT_DDC_DECIMATION : integer := 5;
    constant INT_AVG_MAX_AVERAGE_BY : integer := 5;
    constant INT_MULTIACC_FIFO_DEPTH : integer := 1024;
    constant INT_MULTIACC_CHANNELS : integer := 10;
    constant INT_MULTIACC_REPETITIONS : integer := 15;
    constant INT_CMD_OUTPUT_WIDTH : integer := 5;
    constant INT_MODULE_SELECT_WIDTH : integer := 5;
    constant INT_MODULES_CMD_CNT : integer := 13;
    constant INT_OUT_FIFO_BUFFERS_DEPTH : integer := 1024;

end package generics;



package body generics is 

end package body generics;